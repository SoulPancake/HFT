module VecTest(
  input [0:0] clk
);

  wire [7:0] data_vec[0];
  wire [7:0] data_vec[1];
  wire [7:0] data_vec[2];
  wire [7:0] data_vec[3];

endmodule
