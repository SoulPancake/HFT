module BundleTest(
  input [0:0] clk
);

  wire [7:0] io_bundle_data;
  wire [0:0] io_bundle_valid;

endmodule
