module MemoryTest(
  input [0:0] clk
);

  reg [15:0] data_mem [0:63];

endmodule
