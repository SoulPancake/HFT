module ParameterTest #(
  parameter WIDTH = 8,
  parameter DEPTH = 256
) (
  input [0:0] clk
);

endmodule
