module PolymorphicTest(
);

endmodule
